//
//-------------------------------------------------------------------------------------------------
// filename:  register_file.v
// author:    ikalvarado
// created:   2012-02-20
//-------------------------------------------------------------------------------------------------
// modification history
// author          date        description
// ialvarado       2012-02-20  creation
//-------------------------------------------------------------------------------------------------

//-------------------------------------------------------------------------------------------------
//
// MODULE: register_file
//
//-------------------------------------------------------------------------------------------------
module register_file (
  clock,
  nreset,
  w_en,
  data_in,
  waddr,
  rd_addr_rs,
  rd_addr_rt,
  data_out_rs,
  data_out_rt
);

  //-----------------------------------------------------------------------------------------------
  // Inputs
  //-----------------------------------------------------------------------------------------------
  input clock;
  input nreset;
  input w_en;
  input [04:0] waddr;
  input [04:0] rd_addr_rs;
  input [04:0] rd_addr_rt;
  input [31:0] data_in;

  //-----------------------------------------------------------------------------------------------
  // Outputs
  //-----------------------------------------------------------------------------------------------
  output [31:0] data_out_rs;
  output [31:0] data_out_rt;

  //-----------------------------------------------------------------------------------------------
  // Memory
  //-----------------------------------------------------------------------------------------------
  reg [31:0] memory_array [0:31];
  integer i;

  //-----------------------------------------------------------------------------------------------
  // logic
  //-----------------------------------------------------------------------------------------------
  assign data_out_rs = rd_addr_rs == 0 ? 0 : memory_array[rd_addr_rs];
  assign data_out_rt = rd_addr_rs == 0 ? 0 : memory_array[rd_addr_rt];

  //-----------------------------------------------------------------------------------------------
  // Registers logic
  //-----------------------------------------------------------------------------------------------
  always @(posedge clock, negedge nreset) begin
    if(!nreset) begin
      for(i = 0; i < 32; i = i + 1) begin
        memory_array[i] <= i;
      end
    end
    else begin
      if(w_en) begin
        memory_array[waddr] <= data_in;
      end
    end
  end

endmodule
