//
//-------------------------------------------------------------------------------------------------
// filename:  tag_fifo_optimized.v
// author:    Diana Garcia
// created:   2012-02-26
//-------------------------------------------------------------------------------------------------
// modification history
// author          date        description
// ialvarado       2012-02-26  creation
//-------------------------------------------------------------------------------------------------

//-------------------------------------------------------------------------------------------------
//
// MODULE: tag_fifo_optimized
//
//-------------------------------------------------------------------------------------------------
module tag_fifo_optimized(
  clock,
  nreset,
  flush_valid,
  rd_en,
  wr_en,
  tag_in,
  tag_out,
  tag_fifo_empty
);

  //-----------------------------------------------------------------------------------------------
  // Inputs
  //-----------------------------------------------------------------------------------------------
  input        clock;
  input        nreset;
  input        flush_valid;
  input        rd_en;
  input        wr_en;
  input [04:0] tag_in;

  //-----------------------------------------------------------------------------------------------
  // Outputs
  //-----------------------------------------------------------------------------------------------
  output wire        tag_fifo_empty;
  output wire [04:0] tag_out;

  //-----------------------------------------------------------------------------------------------
  // Internals
  //-----------------------------------------------------------------------------------------------
  reg  [05:0] wp;
  reg  [05:0] rp;
  wire full;

  integer i;
  genvar  n;

  //-----------------------------------------------------------------------------------------------
  // Memory
  //-----------------------------------------------------------------------------------------------
  wire [4:0] memory[0:31];

  assign tag_out        = memory[rp[4:0]];
  assign tag_fifo_empty = wp == rp;
  assign full           = (wp[5] != rp[5]) && wp[4:0] == rp[4:0];

  //-----------------------------------------------------------------------------------------------
  // Memory
  //-----------------------------------------------------------------------------------------------
  generate
    for(n = 0; n < 32; n = n + 1) begin
      assign memory[n] = n[4:0];
    end
  endgenerate

  //-----------------------------------------------------------------------------------------------
  //------ Write Pointer - wp ---------------------------
  //-----------------------------------------------------------------------------------------------
  always @ (posedge clock, negedge nreset) begin
    if(!nreset) begin
      wp <= 32;
    end
    else if(flush_valid) begin
      wp <= 32;
    end
    else begin
      if(wr_en && !full) begin
        wp <= wp + 1;
      end
    end
  end

  //-----------------------------------------------------------------------------------------------
  // ----- Read Pointer - rp ----------------------------
  //-----------------------------------------------------------------------------------------------
  always @ (posedge clock, negedge nreset) begin
    if(!nreset) begin
      rp <= 0;
    end
    else if(flush_valid) begin
      rp <= 0;
    end
    else begin
      if(rd_en && !tag_fifo_empty) begin
        rp <= rp + 1;
      end
    end
  end

endmodule












