
module sync_rom (clock, address, data_out);
  input          clock;
  input  [  4:0] address;
  output [127:0] data_out;

  reg    [127:0] data_out;

  always @(posedge clock) begin
    case (address)
      5'h00:   data_out = 128'h0000002000bf10190080f82000000020;
      5'h01:   data_out = 128'h10c0000c0082302a007f202000001820;
      5'h02:   data_out = 128'h10c0000201cd302a8c8e00008c6d0000;
      5'h03:   data_out = 128'h009f2020007f1820ac8d0000ac6e0000;
      5'h04:   data_out = 128'h08000004005f102210c1fff60082302a;
      5'h05:   data_out = 128'h00bfe019035fd8200000d02000000020;
      5'h06:   data_out = 128'h03ddc82a8f7e00008f5d0000039ae020;
      5'h07:   data_out = 128'h037fd820035fd0201000ffff13200001;
      5'h08:   data_out = 128'h00000020000000201000fff7137c0001;
      5'h09:   data_out = 128'h0121502000bf482000a0102000000020;
      5'h0a:   data_out = 128'h007f68190061202000a0182000003020;
      5'h0b:   data_out = 128'h009f701902e0b02001a060208db70000;
      5'h0c:   data_out = 128'h01c0602010c000020316302a8dd80000;
      5'h0d:   data_out = 128'h1000fff7108a0001008120200300b020;
      5'h0e:   data_out = 128'h00611820ad970000adb6000000000020;
      5'h0f:   data_out = 128'h000000201000ffec1069000100612020;
      5'h10:   data_out = 128'h00bfe019035fd82000bfd01900000020;
      5'h11:   data_out = 128'h03bec82a8f7e00008f5d0000039ae020;
      5'h12:   data_out = 128'h037fd820035fd0201000ffff13390001;
      5'h13:   data_out = 128'h1000ffff000000201000fff7137c0001;
      5'h14:   data_out = 128'h00000020000000200000002000000020;
      5'h15:   data_out = 128'h00000020000000200000002000000020;
      5'h16:   data_out = 128'h00000020000000200000002000000020;
      5'h17:   data_out = 128'h00000020000000200000002000000020;
      5'h18:   data_out = 128'h00000020000000200000002000000020;
      5'h19:   data_out = 128'h00000020000000200000002000000020;
      5'h1a:   data_out = 128'h00000020000000200000002000000020;
      5'h1b:   data_out = 128'h00000020000000200000002000000020;
      5'h1c:   data_out = 128'h00000020000000200000002000000020;
      5'h1d:   data_out = 128'h00000020000000200000002000000020;
      5'h1e:   data_out = 128'h00000020000000200000002000000020;
      5'h1f:   data_out = 128'h00000020000000200000002000000020;
      default: data_out = 128'h1000ffff1000ffff1000ffff1000ffff;
    endcase
  end
endmodule





