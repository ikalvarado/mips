//
//-------------------------------------------------------------------------------------------------
// filename:  i_cache.v
// author:    ikalvarado
// created:   2012-02-03
//-------------------------------------------------------------------------------------------------
// modification history
// author          date        description
// ialvarado       2012-02-03  creation
//-------------------------------------------------------------------------------------------------

//-------------------------------------------------------------------------------------------------
//
// MODULE: i_cache
//
//-------------------------------------------------------------------------------------------------
module i_cache (
  clock,
  nreset,
  rd_en,
  pc_in,
  dout_valid,
  dout
);

  //-----------------------------------------------------------------------------------------------
  // Inputs
  //-----------------------------------------------------------------------------------------------
  input clock;
  input nreset;
  input rd_en;
  input [31:0] pc_in;

  //-----------------------------------------------------------------------------------------------
  // Outputs
  //-----------------------------------------------------------------------------------------------
  output wire dout_valid;
  output wire [127:0] dout;

  //-----------------------------------------------------------------------------------------------
  // Variables
  //-----------------------------------------------------------------------------------------------
  reg         valid_data;

  //-----------------------------------------------------------------------------------------------
  // Initial conditions
  //-----------------------------------------------------------------------------------------------
  sync_rom rom(
    .clock    (clock),
    .address  (pc_in[8:4]),
    .data_out (dout)
  );

  //-----------------------------------------------------------------------------------------------
  // Acknowledge
  //-----------------------------------------------------------------------------------------------
  assign dout_valid = valid_data & rd_en;

  always @(posedge clock) begin
    if(!nreset) begin
      valid_data <= 0;
    end
    else begin
      valid_data <= rd_en;
    end
  end

endmodule
