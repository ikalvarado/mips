//
//-------------------------------------------------------------------------------------------------
// filename:  multiplier_wrapper.v
// author:    lgonzale
// created:   2012-04-05
//-------------------------------------------------------------------------------------------------
// modification history
// author          date        description
// lgonzale        2012-04-06  creation
//-------------------------------------------------------------------------------------------------

//-------------------------------------------------------------------------------------------------
//
// MODULE: multiplier_wrapper
//
//-------------------------------------------------------------------------------------------------
module multiplier_wrapper(
  clock,
  op1,
  op2,
  tag_in,
  out,
  tag_out
);

  //-----------------------------------------------------------------------------------------------
  // input
  //-----------------------------------------------------------------------------------------------
  input        clock;
  input [31:0] op1;
  input [31:0] op2;
  input [ 4:0] tag_in;

  //-----------------------------------------------------------------------------------------------
  // outputs
  //-----------------------------------------------------------------------------------------------
  output wire [31:0] out;
  output wire [ 4:0] tag_out;

  //-----------------------------------------------------------------------------------------------
  // variables
  //-----------------------------------------------------------------------------------------------
  reg  [ 4:0] tag_st[ 2:0];
  integer i;
  
  assign tag_out = tag_st[2];
  
  signed_multiplier core_multiplier(
    .out( out       ),
    .clk( clock     ),
    .a  ( op1[15:0] ),
    .b  ( op2[15:0] )
  );

  //-----------------------------------------------------------------------------------------------
  // logic
  //-----------------------------------------------------------------------------------------------
  always @(posedge clock)  begin
    tag_st[0] <= tag_in;
    for(i = 1; i < 3; i = i + 1) begin
      tag_st[i] <= tag_st[i - 1];
    end
  end

endmodule



